`include "../common/structs/core_structures.sv"

module tych_ing (

input wire clk,
input wire reset,

input wire core_avl_t core_avl_in [1:0],
output core_avl_t core_avl_out [1:0]
);


endmodule