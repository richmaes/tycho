module tych_ing

input logic clk,
input logic reset,

input core_avl_t core_avl_in [1:0],
output core_avl_t core_avl_out [1:0]
);


endmodule