module tych_egr (
input logic clk,
input logic reset
);

endmodule